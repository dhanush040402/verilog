module AND_2(output Y, input A, B);
    and(Y, A, B); 
endmodule
